// $Id: $mg68
// File name:   tb_discrimination_parameter_creator.sv
// Created:     23/11/2014
// Author:      Tatsu
// Lab Section: 337-02
// Version:     1.0  Initial Design Entry
// Description: Finds the discrimination parameter!

`timescale 1ns / 100ps // Time unit of one nanosecond, with a precision of 100ps.

module tb_discrimination_parameter_creator();

	parameter CLK_PERIOD = 10; // 100 MHz input.

	// Inputs as registers.
	reg tb_clk;
	reg tb_nrst;
	reg [19:0] tb_data_input;
	reg [19:0] tb_baseline_value;
	
	// Outputs as wires.
	wire [25:0] tb_discrimination_parameter;
	
	discrimination_parameter_creator Dd 
	(
		.clk (tb_clk),
		.nrst (tb_nrst),
	 	.data_input (tb_data_input),
	 	.baseline_value (tb_baseline_value),
	 	.discrimination_parameter (tb_discrimination_parameter)
	); // Device Under Test

	always 
	begin : CLOCK_GENERATION
		tb_clk = 1'b0;
		#(CLK_PERIOD / 2); // 5ns
		tb_clk = 1'b1;
		#(CLK_PERIOD / 2); // 5ns
	end

	initial // Testbench time!
	begin : TESTING_THE_DISCRIMINATOR // "I'll be back!"

		assign tb_nrst = 1'b1; // Default value.
		assign tb_data_input = 0; // Default value.
		assign tb_baseline_value = 0; // Default value.

		#(2 * CLK_PERIOD); // Get away from time = 0.

		assign tb_nrst = 1'b0; // Reset!

		#(2 * CLK_PERIOD);

		assign tb_nrst = 1'b1; // Default value.

		/* === Test Case 1 === */

		assign tb_data_input = 21300;
		assign tb_baseline_value = 12500;

		#(CLK_PERIOD);

		assign tb_data_input = 21301;
		#(CLK_PERIOD);
		assign tb_data_input = 21302;
		#(CLK_PERIOD);
		assign tb_data_input = 21303;
		#(CLK_PERIOD);
		assign tb_data_input = 21304;
		#(CLK_PERIOD);
		assign tb_data_input = 21305;
		#(CLK_PERIOD);
		assign tb_data_input = 21306;
		#(CLK_PERIOD);
		assign tb_data_input = 21307;
		#(CLK_PERIOD);
		assign tb_data_input = 21308;
		#(CLK_PERIOD);
		assign tb_data_input = 21309;
		#(CLK_PERIOD);
		assign tb_data_input = 21310;
		#(CLK_PERIOD);
		assign tb_data_input = 21311;
		#(CLK_PERIOD);
		assign tb_data_input = 21312;
		#(CLK_PERIOD);
		assign tb_data_input = 21313;
		#(CLK_PERIOD);
		assign tb_data_input = 21314;
		#(CLK_PERIOD);
		assign tb_data_input = 21315;
		#(CLK_PERIOD);
		assign tb_data_input = 21316;
		#(CLK_PERIOD);
		assign tb_data_input = 21317;
		#(CLK_PERIOD);
		assign tb_data_input = 21318;
		#(CLK_PERIOD);
		assign tb_data_input = 21319;
		#(CLK_PERIOD);
		assign tb_data_input = 21320;
		#(CLK_PERIOD);
		assign tb_data_input = 21321;
		#(CLK_PERIOD);
		assign tb_data_input = 21322;
		#(CLK_PERIOD);
		assign tb_data_input = 21323;
		#(CLK_PERIOD);
		assign tb_data_input = 21324;
		#(CLK_PERIOD);
		assign tb_data_input = 21325;
		#(CLK_PERIOD);
		assign tb_data_input = 21326;
		#(CLK_PERIOD);
		assign tb_data_input = 21327;
		#(CLK_PERIOD);
		assign tb_data_input = 21328;
		#(CLK_PERIOD);
		assign tb_data_input = 21329;
		#(CLK_PERIOD);
		assign tb_data_input = 21330;
		#(CLK_PERIOD);
		assign tb_data_input = 21331;
		#(CLK_PERIOD);
		assign tb_data_input = 21332;
		#(CLK_PERIOD);
		assign tb_data_input = 21333;
		#(CLK_PERIOD);
		assign tb_data_input = 21334;
		#(CLK_PERIOD);
		assign tb_data_input = 21335;
		#(CLK_PERIOD);
		assign tb_data_input = 21336;
		#(CLK_PERIOD);
		assign tb_data_input = 21337;
		#(CLK_PERIOD);
		assign tb_data_input = 21338;
		#(CLK_PERIOD);
		assign tb_data_input = 21339;
		#(CLK_PERIOD);
		assign tb_data_input = 21340;
		#(CLK_PERIOD);
		assign tb_data_input = 21341;
		#(CLK_PERIOD);
		assign tb_data_input = 21342;
		#(CLK_PERIOD);
		assign tb_data_input = 21343;
		#(CLK_PERIOD);
		assign tb_data_input = 21344;
		#(CLK_PERIOD);
		assign tb_data_input = 21345;
		#(CLK_PERIOD);
		assign tb_data_input = 21346;
		#(CLK_PERIOD);
		assign tb_data_input = 21347;
		#(CLK_PERIOD);
		assign tb_data_input = 21348;
		#(CLK_PERIOD);
		assign tb_data_input = 21349;
		#(CLK_PERIOD);
		assign tb_data_input = 21350;
		#(CLK_PERIOD);
		assign tb_data_input = 21351;
		#(CLK_PERIOD);
		assign tb_data_input = 21352;
		#(CLK_PERIOD);
		assign tb_data_input = 21353;
		#(CLK_PERIOD);
		assign tb_data_input = 21354;
		#(CLK_PERIOD);
		assign tb_data_input = 21355;
		#(CLK_PERIOD);
		assign tb_data_input = 21356;
		#(CLK_PERIOD);
		assign tb_data_input = 21357;
		#(CLK_PERIOD);
		assign tb_data_input = 21358;
		#(CLK_PERIOD);
		assign tb_data_input = 21359;
		#(CLK_PERIOD);
		assign tb_data_input = 21360;
		#(CLK_PERIOD);
		assign tb_data_input = 21361;
		#(CLK_PERIOD);
		assign tb_data_input = 21362;
		#(CLK_PERIOD);
		assign tb_data_input = 21363;
		#(CLK_PERIOD);
		assign tb_data_input = 21364;
		#(CLK_PERIOD);
		assign tb_data_input = 21365;
		#(CLK_PERIOD);
		assign tb_data_input = 21366;
		#(CLK_PERIOD);
		assign tb_data_input = 21367;
		#(CLK_PERIOD);
		assign tb_data_input = 21368;
		#(CLK_PERIOD);
		assign tb_data_input = 21369;
		#(CLK_PERIOD);
		assign tb_data_input = 21370;
		#(CLK_PERIOD);
		assign tb_data_input = 21371;
		#(CLK_PERIOD);
		assign tb_data_input = 21372;
		#(CLK_PERIOD);
		assign tb_data_input = 21373;
		#(CLK_PERIOD);
		assign tb_data_input = 21374;
		#(CLK_PERIOD);
		assign tb_data_input = 21375;
		#(CLK_PERIOD);
		assign tb_data_input = 21376;
		#(CLK_PERIOD);
		assign tb_data_input = 21377;
		#(CLK_PERIOD);
		assign tb_data_input = 21378;
		#(CLK_PERIOD);
		assign tb_data_input = 21379;
		#(CLK_PERIOD);
		assign tb_data_input = 21380;
		#(CLK_PERIOD);
		assign tb_data_input = 21381;
		#(CLK_PERIOD);
		assign tb_data_input = 21382;
		#(CLK_PERIOD);
		assign tb_data_input = 21383;
		#(CLK_PERIOD);
		assign tb_data_input = 21384;
		#(CLK_PERIOD);
		assign tb_data_input = 21385;
		#(CLK_PERIOD);
		assign tb_data_input = 21386;
		#(CLK_PERIOD);
		assign tb_data_input = 21387;
		#(CLK_PERIOD);
		assign tb_data_input = 21388;
		#(CLK_PERIOD);
		assign tb_data_input = 21389;
		#(CLK_PERIOD);
		assign tb_data_input = 21390;
		#(CLK_PERIOD);
		assign tb_data_input = 21391;
		#(CLK_PERIOD);
		assign tb_data_input = 21392;
		#(CLK_PERIOD);
		assign tb_data_input = 21393;
		#(CLK_PERIOD);
		assign tb_data_input = 21394;
		#(CLK_PERIOD);
		assign tb_data_input = 21395;
		#(CLK_PERIOD);
		assign tb_data_input = 21396;
		#(CLK_PERIOD);
		assign tb_data_input = 21397;
		#(CLK_PERIOD);
		assign tb_data_input = 21398;
		#(CLK_PERIOD);
		assign tb_data_input = 21399;
		#(CLK_PERIOD);
		assign tb_data_input = 21400;
		#(CLK_PERIOD);
		assign tb_data_input = 21401;
		#(CLK_PERIOD);
		assign tb_data_input = 21402;
		#(CLK_PERIOD);
		assign tb_data_input = 21403;
		#(CLK_PERIOD);
		assign tb_data_input = 21404;
		#(CLK_PERIOD);
		assign tb_data_input = 21405;
		#(CLK_PERIOD);
		assign tb_data_input = 21406;
		#(CLK_PERIOD);
		assign tb_data_input = 21407;
		#(CLK_PERIOD);
		assign tb_data_input = 21408;
		#(CLK_PERIOD);
		assign tb_data_input = 21409;
		#(CLK_PERIOD);
		assign tb_data_input = 21410;
		#(CLK_PERIOD);
		assign tb_data_input = 21411;
		#(CLK_PERIOD);
		assign tb_data_input = 21412;
		#(CLK_PERIOD);
		assign tb_data_input = 21413;
		#(CLK_PERIOD);
		assign tb_data_input = 21414;
		#(CLK_PERIOD);
		assign tb_data_input = 21415;
		#(CLK_PERIOD);
		assign tb_data_input = 21416;
		#(CLK_PERIOD);
		assign tb_data_input = 21417;
		#(CLK_PERIOD);
		assign tb_data_input = 21418;
		#(CLK_PERIOD);
		assign tb_data_input = 21419;
		#(CLK_PERIOD);
		assign tb_data_input = 21420;
		#(CLK_PERIOD);
		assign tb_data_input = 21421;
		#(CLK_PERIOD);
		assign tb_data_input = 21422;
		#(CLK_PERIOD);
		assign tb_data_input = 21423;
		#(CLK_PERIOD);
		assign tb_data_input = 21424;
		#(CLK_PERIOD);
		assign tb_data_input = 21425;
		#(CLK_PERIOD);
		assign tb_data_input = 21426;
		#(CLK_PERIOD);
		assign tb_data_input = 21427;
		#(CLK_PERIOD);
		assign tb_data_input = 21428;
		#(CLK_PERIOD);
		assign tb_data_input = 21429;
		#(CLK_PERIOD);
		assign tb_data_input = 21430;
		#(CLK_PERIOD);
		assign tb_data_input = 21431;
		#(CLK_PERIOD);
		assign tb_data_input = 21432;
		#(CLK_PERIOD);
		assign tb_data_input = 21433;
		#(CLK_PERIOD);
		assign tb_data_input = 21434;
		#(CLK_PERIOD);
		assign tb_data_input = 21435;
		#(CLK_PERIOD);
		assign tb_data_input = 21436;
		#(CLK_PERIOD);
		assign tb_data_input = 21437;
		#(CLK_PERIOD);
		assign tb_data_input = 21438;
		#(CLK_PERIOD);
		assign tb_data_input = 21439;
		#(CLK_PERIOD);
		assign tb_data_input = 21440;
		#(CLK_PERIOD);
		assign tb_data_input = 21441;
		#(CLK_PERIOD);
		assign tb_data_input = 21442;
		#(CLK_PERIOD);
		assign tb_data_input = 21443;
		#(CLK_PERIOD);
		assign tb_data_input = 21444;
		#(CLK_PERIOD);
		assign tb_data_input = 21445;
		#(CLK_PERIOD);
		assign tb_data_input = 21446;
		#(CLK_PERIOD);
		assign tb_data_input = 21447;
		#(CLK_PERIOD);
		assign tb_data_input = 21448;
		#(CLK_PERIOD);
		assign tb_data_input = 21449;
		#(CLK_PERIOD);
		assign tb_data_input = 21450;
		#(CLK_PERIOD);
		assign tb_data_input = 21451;
		#(CLK_PERIOD);
		assign tb_data_input = 21452;
		#(CLK_PERIOD);
		assign tb_data_input = 21453;
		#(CLK_PERIOD);
		assign tb_data_input = 21454;
		#(CLK_PERIOD);
		assign tb_data_input = 21455;
		#(CLK_PERIOD);
		assign tb_data_input = 21456;
		#(CLK_PERIOD);
		assign tb_data_input = 21457;
		#(CLK_PERIOD);
		assign tb_data_input = 21458;
		#(CLK_PERIOD);
		assign tb_data_input = 21459;
		#(CLK_PERIOD);
		assign tb_data_input = 21460;
		#(CLK_PERIOD);
		assign tb_data_input = 21461;
		#(CLK_PERIOD);
		assign tb_data_input = 21462;
		#(CLK_PERIOD);
		assign tb_data_input = 21463;
		#(CLK_PERIOD);
		assign tb_data_input = 21464;
		#(CLK_PERIOD);
		assign tb_data_input = 21465;
		#(CLK_PERIOD);
		assign tb_data_input = 21466;
		#(CLK_PERIOD);
		assign tb_data_input = 21467;
		#(CLK_PERIOD);
		assign tb_data_input = 21468;
		#(CLK_PERIOD);
		assign tb_data_input = 21469;
		#(CLK_PERIOD);
		assign tb_data_input = 21470;
		#(CLK_PERIOD);
		assign tb_data_input = 21471;
		#(CLK_PERIOD);
		assign tb_data_input = 21472;
		#(CLK_PERIOD);
		assign tb_data_input = 21473;
		#(CLK_PERIOD);
		assign tb_data_input = 21474;
		#(CLK_PERIOD);
		assign tb_data_input = 21475;
		#(CLK_PERIOD);
		assign tb_data_input = 21476;
		#(CLK_PERIOD);
		assign tb_data_input = 21477;
		#(CLK_PERIOD);
		assign tb_data_input = 21478;
		#(CLK_PERIOD);
		assign tb_data_input = 21479;
		#(CLK_PERIOD);
		assign tb_data_input = 21480;
		#(CLK_PERIOD);
		assign tb_data_input = 21481;
		#(CLK_PERIOD);
		assign tb_data_input = 21482;
		#(CLK_PERIOD);
		assign tb_data_input = 21483;
		#(CLK_PERIOD);
		assign tb_data_input = 21484;
		#(CLK_PERIOD);
		assign tb_data_input = 21485;
		#(CLK_PERIOD);
		assign tb_data_input = 21486;
		#(CLK_PERIOD);
		assign tb_data_input = 21487;
		#(CLK_PERIOD);
		assign tb_data_input = 21488;
		#(CLK_PERIOD);
		assign tb_data_input = 21489;
		#(CLK_PERIOD);
		assign tb_data_input = 21490;
		#(CLK_PERIOD);
		assign tb_data_input = 21491;
		#(CLK_PERIOD);
		assign tb_data_input = 21492;
		#(CLK_PERIOD);
		assign tb_data_input = 21493;
		#(CLK_PERIOD);
		assign tb_data_input = 21494;
		#(CLK_PERIOD);
		assign tb_data_input = 21495;
		#(CLK_PERIOD);
		assign tb_data_input = 21496;
		#(CLK_PERIOD);
		assign tb_data_input = 21497;
		#(CLK_PERIOD);
		assign tb_data_input = 21498;
		#(CLK_PERIOD);
		assign tb_data_input = 21499;
		#(CLK_PERIOD);
		assign tb_data_input = 21500;
		#(CLK_PERIOD);
		assign tb_data_input = 21501;
		#(CLK_PERIOD);
		assign tb_data_input = 21502;
		#(CLK_PERIOD);
		assign tb_data_input = 21503;
		#(CLK_PERIOD);
		assign tb_data_input = 21504;
		#(CLK_PERIOD);
		assign tb_data_input = 21505;
		#(CLK_PERIOD);
		assign tb_data_input = 21506;
		#(CLK_PERIOD);
		assign tb_data_input = 21507;
		#(CLK_PERIOD);
		assign tb_data_input = 21508;
		#(CLK_PERIOD);
		assign tb_data_input = 21509;
		#(CLK_PERIOD);
		assign tb_data_input = 21510;
		#(CLK_PERIOD);
		assign tb_data_input = 21511;
		#(CLK_PERIOD);
		assign tb_data_input = 21512;
		#(CLK_PERIOD);
		assign tb_data_input = 21513;
		#(CLK_PERIOD);
		assign tb_data_input = 21514;
		#(CLK_PERIOD);
		assign tb_data_input = 21515;
		#(CLK_PERIOD);
		assign tb_data_input = 21516;
		#(CLK_PERIOD);
		assign tb_data_input = 21517;
		#(CLK_PERIOD);
		assign tb_data_input = 21518;
		#(CLK_PERIOD);
		assign tb_data_input = 21519;
		#(CLK_PERIOD);
		assign tb_data_input = 21520;
		#(CLK_PERIOD);
		assign tb_data_input = 21521;
		#(CLK_PERIOD);
		assign tb_data_input = 21522;
		#(CLK_PERIOD);
		assign tb_data_input = 21523;
		#(CLK_PERIOD);
		assign tb_data_input = 21524;
		#(CLK_PERIOD);
		assign tb_data_input = 21525;
		#(CLK_PERIOD);
		assign tb_data_input = 21526;
		#(CLK_PERIOD);
		assign tb_data_input = 21527;
		#(CLK_PERIOD);
		assign tb_data_input = 21528;
		#(CLK_PERIOD);
		assign tb_data_input = 21529;
		#(CLK_PERIOD);
		assign tb_data_input = 21530;
		#(CLK_PERIOD);
		assign tb_data_input = 21531;
		#(CLK_PERIOD);
		assign tb_data_input = 21532;
		#(CLK_PERIOD);
		assign tb_data_input = 21533;
		#(CLK_PERIOD);
		assign tb_data_input = 21534;
		#(CLK_PERIOD);
		assign tb_data_input = 21535;
		#(CLK_PERIOD);
		assign tb_data_input = 21536;
		#(CLK_PERIOD);
		assign tb_data_input = 21537;
		#(CLK_PERIOD);
		assign tb_data_input = 21538;
		#(CLK_PERIOD);
		assign tb_data_input = 21539;
		#(CLK_PERIOD);
		assign tb_data_input = 21540;
		#(CLK_PERIOD);
		assign tb_data_input = 21541;
		#(CLK_PERIOD);
		assign tb_data_input = 21542;
		#(CLK_PERIOD);
		assign tb_data_input = 21543;
		#(CLK_PERIOD);
		assign tb_data_input = 21544;
		#(CLK_PERIOD);
		assign tb_data_input = 21545;
		#(CLK_PERIOD);
		assign tb_data_input = 21546;
		#(CLK_PERIOD);
		assign tb_data_input = 21547;
		#(CLK_PERIOD);
		assign tb_data_input = 21548;
		#(CLK_PERIOD);
		assign tb_data_input = 21549;
		#(CLK_PERIOD);
		assign tb_data_input = 21550;
		#(CLK_PERIOD);
		assign tb_data_input = 21551;
		#(CLK_PERIOD);
		assign tb_data_input = 21552;
		#(CLK_PERIOD);
		assign tb_data_input = 21553;
		#(CLK_PERIOD);
		assign tb_data_input = 21554;
		#(CLK_PERIOD);
		assign tb_data_input = 21555;
		#(CLK_PERIOD);
		assign tb_data_input = 21556;
		#(CLK_PERIOD);
		assign tb_data_input = 21557;
		#(CLK_PERIOD);
		assign tb_data_input = 21558;
		#(CLK_PERIOD);
		assign tb_data_input = 21559;
		#(CLK_PERIOD);
		assign tb_data_input = 21560;
		#(CLK_PERIOD);
		assign tb_data_input = 21561;
		#(CLK_PERIOD);
		assign tb_data_input = 21562;
		#(CLK_PERIOD);
		assign tb_data_input = 21563;
		#(CLK_PERIOD);
		assign tb_data_input = 21564;
		#(CLK_PERIOD);
		assign tb_data_input = 21565;
		#(CLK_PERIOD);
		assign tb_data_input = 21566;
		#(CLK_PERIOD);
		assign tb_data_input = 21567;
		#(CLK_PERIOD);
		assign tb_data_input = 21568;
		#(CLK_PERIOD);
		assign tb_data_input = 21569;
		#(CLK_PERIOD);
		assign tb_data_input = 21570;
		#(CLK_PERIOD);
		assign tb_data_input = 21571;
		#(CLK_PERIOD);
		assign tb_data_input = 21572;
		#(CLK_PERIOD);
		assign tb_data_input = 21573;
		#(CLK_PERIOD);
		assign tb_data_input = 21574;
		#(CLK_PERIOD);
		assign tb_data_input = 21575;
		#(CLK_PERIOD);
		assign tb_data_input = 21576;
		#(CLK_PERIOD);
		assign tb_data_input = 21577;
		#(CLK_PERIOD);
		assign tb_data_input = 21578;
		#(CLK_PERIOD);
		assign tb_data_input = 21579;
		#(CLK_PERIOD);
		assign tb_data_input = 21580;
		#(CLK_PERIOD);
		assign tb_data_input = 21581;
		#(CLK_PERIOD);
		assign tb_data_input = 21582;
		#(CLK_PERIOD);
		assign tb_data_input = 21583;
		#(CLK_PERIOD);
		assign tb_data_input = 21584;
		#(CLK_PERIOD);
		assign tb_data_input = 21585;
		#(CLK_PERIOD);
		assign tb_data_input = 21586;
		#(CLK_PERIOD);
		assign tb_data_input = 21587;
		#(CLK_PERIOD);
		assign tb_data_input = 21588;
		#(CLK_PERIOD);
		assign tb_data_input = 21589;
		#(CLK_PERIOD);
		assign tb_data_input = 21590;
		#(CLK_PERIOD);
		assign tb_data_input = 21591;
		#(CLK_PERIOD);
		assign tb_data_input = 21592;
		#(CLK_PERIOD);
		assign tb_data_input = 21593;
		#(CLK_PERIOD);
		assign tb_data_input = 21594;
		#(CLK_PERIOD);
		assign tb_data_input = 21595;
		#(CLK_PERIOD);
		assign tb_data_input = 21596;
		#(CLK_PERIOD);
		assign tb_data_input = 21597;
		#(CLK_PERIOD);
		assign tb_data_input = 21598;
		#(CLK_PERIOD);
		assign tb_data_input = 21599;
		#(CLK_PERIOD);
		assign tb_data_input = 21600;
		#(CLK_PERIOD);
		assign tb_data_input = 21601;
		#(CLK_PERIOD);
		assign tb_data_input = 21602;
		#(CLK_PERIOD);
		assign tb_data_input = 21603;
		#(CLK_PERIOD);
		assign tb_data_input = 21604;
		#(CLK_PERIOD);
		assign tb_data_input = 21605;
		#(CLK_PERIOD);
		assign tb_data_input = 21606;
		#(CLK_PERIOD);
		assign tb_data_input = 21607;
		#(CLK_PERIOD);
		assign tb_data_input = 21608;
		#(CLK_PERIOD);
		assign tb_data_input = 21609;
		#(CLK_PERIOD);
		assign tb_data_input = 21610;
		#(CLK_PERIOD);
		assign tb_data_input = 21611;
		#(CLK_PERIOD);
		assign tb_data_input = 21612;
		#(CLK_PERIOD);
		assign tb_data_input = 21613;
		#(CLK_PERIOD);
		assign tb_data_input = 21614;
		#(CLK_PERIOD);
		assign tb_data_input = 21615;
		#(CLK_PERIOD);
		assign tb_data_input = 21616;
		#(CLK_PERIOD);
		assign tb_data_input = 21617;
		#(CLK_PERIOD);
		assign tb_data_input = 21618;
		#(CLK_PERIOD);
		assign tb_data_input = 21619;
		#(CLK_PERIOD);
		assign tb_data_input = 21620;
		#(CLK_PERIOD);
		assign tb_data_input = 21621;
		#(CLK_PERIOD);
		assign tb_data_input = 21622;
		#(CLK_PERIOD);
		assign tb_data_input = 21623;
		#(CLK_PERIOD);
		assign tb_data_input = 21624;
		#(CLK_PERIOD);
		assign tb_data_input = 21625;
		#(CLK_PERIOD);
		assign tb_data_input = 21626;
		#(CLK_PERIOD);
		assign tb_data_input = 21627;
		#(CLK_PERIOD);
		assign tb_data_input = 21628;
		#(CLK_PERIOD);
		assign tb_data_input = 21629;
		#(CLK_PERIOD);
		assign tb_data_input = 21630;
		#(CLK_PERIOD);
		assign tb_data_input = 21631;
		#(CLK_PERIOD);
		assign tb_data_input = 21632;
		#(CLK_PERIOD);
		assign tb_data_input = 21633;
		#(CLK_PERIOD);
		assign tb_data_input = 21634;
		#(CLK_PERIOD);
		assign tb_data_input = 21635;
		#(CLK_PERIOD);
		assign tb_data_input = 21636;
		#(CLK_PERIOD);
		assign tb_data_input = 21637;
		#(CLK_PERIOD);
		assign tb_data_input = 21638;
		#(CLK_PERIOD);
		assign tb_data_input = 21639;
		#(CLK_PERIOD);
		assign tb_data_input = 21640;
		#(CLK_PERIOD);
		assign tb_data_input = 21641;
		#(CLK_PERIOD);
		assign tb_data_input = 21642;
		#(CLK_PERIOD);
		assign tb_data_input = 21643;
		#(CLK_PERIOD);
		assign tb_data_input = 21644;
		#(CLK_PERIOD);
		assign tb_data_input = 21645;
		#(CLK_PERIOD);
		assign tb_data_input = 21646;
		#(CLK_PERIOD);
		assign tb_data_input = 21647;
		#(CLK_PERIOD);
		assign tb_data_input = 21648;
		#(CLK_PERIOD);
		assign tb_data_input = 21649;
		#(CLK_PERIOD);
		assign tb_data_input = 21650;
		#(CLK_PERIOD);
		assign tb_data_input = 21651;
		#(CLK_PERIOD);
		assign tb_data_input = 21652;
		#(CLK_PERIOD);
		assign tb_data_input = 21653;
		#(CLK_PERIOD);
		assign tb_data_input = 21654;
		#(CLK_PERIOD);
		assign tb_data_input = 21655;
		#(CLK_PERIOD);
		assign tb_data_input = 21656;
		#(CLK_PERIOD);
		assign tb_data_input = 21657;
		#(CLK_PERIOD);
		assign tb_data_input = 21658;
		#(CLK_PERIOD);
		assign tb_data_input = 21659;
		#(CLK_PERIOD);
		assign tb_data_input = 21660;
		#(CLK_PERIOD);
		assign tb_data_input = 21661;
		#(CLK_PERIOD);
		assign tb_data_input = 21662;
		#(CLK_PERIOD);
		assign tb_data_input = 21663;
		#(CLK_PERIOD);
		assign tb_data_input = 21664;
		#(CLK_PERIOD);
		assign tb_data_input = 21665;
		#(CLK_PERIOD);
		assign tb_data_input = 21666;
		#(CLK_PERIOD);
		assign tb_data_input = 21667;
		#(CLK_PERIOD);
		assign tb_data_input = 21668;
		#(CLK_PERIOD);
		assign tb_data_input = 21669;
		#(CLK_PERIOD);
		assign tb_data_input = 21670;
		#(CLK_PERIOD);
		assign tb_data_input = 21671;
		#(CLK_PERIOD);
		assign tb_data_input = 21672;
		#(CLK_PERIOD);
		assign tb_data_input = 21673;
		#(CLK_PERIOD);
		assign tb_data_input = 21674;
		#(CLK_PERIOD);
		assign tb_data_input = 21675;
		#(CLK_PERIOD);
		assign tb_data_input = 21676;
		#(CLK_PERIOD);
		assign tb_data_input = 21677;
		#(CLK_PERIOD);
		assign tb_data_input = 21678;
		#(CLK_PERIOD);
		assign tb_data_input = 21679;
		#(CLK_PERIOD);
		assign tb_data_input = 21680;
		#(CLK_PERIOD);
		assign tb_data_input = 21681;
		#(CLK_PERIOD);
		assign tb_data_input = 21682;
		#(CLK_PERIOD);
		assign tb_data_input = 21683;
		#(CLK_PERIOD);
		assign tb_data_input = 21684;
		#(CLK_PERIOD);
		assign tb_data_input = 21685;
		#(CLK_PERIOD);
		assign tb_data_input = 21686;
		#(CLK_PERIOD);
		assign tb_data_input = 21687;
		#(CLK_PERIOD);
		assign tb_data_input = 21688;
		#(CLK_PERIOD);
		assign tb_data_input = 21689;
		#(CLK_PERIOD);
		assign tb_data_input = 21690;
		#(CLK_PERIOD);
		assign tb_data_input = 21691;
		#(CLK_PERIOD);
		assign tb_data_input = 21692;
		#(CLK_PERIOD);
		assign tb_data_input = 21693;
		#(CLK_PERIOD);
		assign tb_data_input = 21694;
		#(CLK_PERIOD);
		assign tb_data_input = 21695;
		#(CLK_PERIOD);
		assign tb_data_input = 21696;
		#(CLK_PERIOD);
		assign tb_data_input = 21697;
		#(CLK_PERIOD);
		assign tb_data_input = 21698;
		#(CLK_PERIOD);
		assign tb_data_input = 21699;
		#(CLK_PERIOD);
		assign tb_data_input = 21700;
		#(CLK_PERIOD);
		assign tb_data_input = 21701;
		#(CLK_PERIOD);
		assign tb_data_input = 21702;
		#(CLK_PERIOD);
		assign tb_data_input = 21703;
		#(CLK_PERIOD);
		assign tb_data_input = 21704;
		#(CLK_PERIOD);
		assign tb_data_input = 21705;
		#(CLK_PERIOD);
		assign tb_data_input = 21706;
		#(CLK_PERIOD);
		assign tb_data_input = 21707;
		#(CLK_PERIOD);
		assign tb_data_input = 21708;
		#(CLK_PERIOD);
		assign tb_data_input = 21709;
		#(CLK_PERIOD);
		assign tb_data_input = 21710;
		#(CLK_PERIOD);
		assign tb_data_input = 21711;
		#(CLK_PERIOD);
		assign tb_data_input = 21712;
		#(CLK_PERIOD);
		assign tb_data_input = 21713;
		#(CLK_PERIOD);
		assign tb_data_input = 21714;
		#(CLK_PERIOD);
		assign tb_data_input = 21715;
		#(CLK_PERIOD);
		assign tb_data_input = 21716;
		#(CLK_PERIOD);
		assign tb_data_input = 21717;
		#(CLK_PERIOD);
		assign tb_data_input = 21718;
		#(CLK_PERIOD);
		assign tb_data_input = 21719;
		#(CLK_PERIOD);
		assign tb_data_input = 21720;
		#(CLK_PERIOD);
		assign tb_data_input = 21721;
		#(CLK_PERIOD);
		assign tb_data_input = 21722;
		#(CLK_PERIOD);
		assign tb_data_input = 21723;
		#(CLK_PERIOD);
		assign tb_data_input = 21724;
		#(CLK_PERIOD);
		assign tb_data_input = 21725;
		#(CLK_PERIOD);
		assign tb_data_input = 21726;
		#(CLK_PERIOD);
		assign tb_data_input = 21727;
		#(CLK_PERIOD);
		assign tb_data_input = 21728;
		#(CLK_PERIOD);
		assign tb_data_input = 21729;
		#(CLK_PERIOD);
		assign tb_data_input = 21730;
		#(CLK_PERIOD);
		assign tb_data_input = 21731;
		#(CLK_PERIOD);
		assign tb_data_input = 21732;
		#(CLK_PERIOD);
		assign tb_data_input = 21733;
		#(CLK_PERIOD);
		assign tb_data_input = 21734;
		#(CLK_PERIOD);
		assign tb_data_input = 21735;
		#(CLK_PERIOD);
		assign tb_data_input = 21736;
		#(CLK_PERIOD);
		assign tb_data_input = 21737;
		#(CLK_PERIOD);
		assign tb_data_input = 21738;
		#(CLK_PERIOD);
		assign tb_data_input = 21739;
		#(CLK_PERIOD);
		assign tb_data_input = 21740;
		#(CLK_PERIOD);
		assign tb_data_input = 21741;
		#(CLK_PERIOD);
		assign tb_data_input = 21742;
		#(CLK_PERIOD);
		assign tb_data_input = 21743;
		#(CLK_PERIOD);
		assign tb_data_input = 21744;
		#(CLK_PERIOD);
		assign tb_data_input = 21745;
		#(CLK_PERIOD);
		assign tb_data_input = 21746;
		#(CLK_PERIOD);
		assign tb_data_input = 21747;
		#(CLK_PERIOD);
		assign tb_data_input = 21748;
		#(CLK_PERIOD);
		assign tb_data_input = 21749;
		#(CLK_PERIOD);
		assign tb_data_input = 21750;
		#(CLK_PERIOD);
		assign tb_data_input = 21751;
		#(CLK_PERIOD);
		assign tb_data_input = 21752;
		#(CLK_PERIOD);
		assign tb_data_input = 21753;
		#(CLK_PERIOD);
		assign tb_data_input = 21754;
		#(CLK_PERIOD);
		assign tb_data_input = 21755;
		#(CLK_PERIOD);
		assign tb_data_input = 21756;
		#(CLK_PERIOD);
		assign tb_data_input = 21757;
		#(CLK_PERIOD);
		assign tb_data_input = 21758;
		#(CLK_PERIOD);
		assign tb_data_input = 21759;
		#(CLK_PERIOD);
		assign tb_data_input = 21760;
		#(CLK_PERIOD);
		assign tb_data_input = 21761;
		#(CLK_PERIOD);
		assign tb_data_input = 21762;
		#(CLK_PERIOD);
		assign tb_data_input = 21763;
		#(CLK_PERIOD);
		assign tb_data_input = 21764;
		#(CLK_PERIOD);
		assign tb_data_input = 21765;
		#(CLK_PERIOD);
		assign tb_data_input = 21766;
		#(CLK_PERIOD);
		assign tb_data_input = 21767;
		#(CLK_PERIOD);
		assign tb_data_input = 21768;
		#(CLK_PERIOD);
		assign tb_data_input = 21769;
		#(CLK_PERIOD);
		assign tb_data_input = 21770;
		#(CLK_PERIOD);
		assign tb_data_input = 21771;
		#(CLK_PERIOD);
		assign tb_data_input = 21772;
		#(CLK_PERIOD);
		assign tb_data_input = 21773;
		#(CLK_PERIOD);
		assign tb_data_input = 21774;
		#(CLK_PERIOD);
		assign tb_data_input = 21775;
		#(CLK_PERIOD);
		assign tb_data_input = 21776;
		#(CLK_PERIOD);
		assign tb_data_input = 21777;
		#(CLK_PERIOD);
		assign tb_data_input = 21778;
		#(CLK_PERIOD);
		assign tb_data_input = 21779;
		#(CLK_PERIOD);
		assign tb_data_input = 21780;
		#(CLK_PERIOD);
		assign tb_data_input = 21781;
		#(CLK_PERIOD);
		assign tb_data_input = 21782;
		#(CLK_PERIOD);
		assign tb_data_input = 21783;
		#(CLK_PERIOD);
		assign tb_data_input = 21784;
		#(CLK_PERIOD);
		assign tb_data_input = 21785;
		#(CLK_PERIOD);
		assign tb_data_input = 21786;
		#(CLK_PERIOD);
		assign tb_data_input = 21787;
		#(CLK_PERIOD);
		assign tb_data_input = 21788;
		#(CLK_PERIOD);
		assign tb_data_input = 21789;
		#(CLK_PERIOD);
		assign tb_data_input = 21790;
		#(CLK_PERIOD);
		assign tb_data_input = 21791;
		#(CLK_PERIOD);
		assign tb_data_input = 21792;
		#(CLK_PERIOD);
		assign tb_data_input = 21793;
		#(CLK_PERIOD);
		assign tb_data_input = 21794;
		#(CLK_PERIOD);
		assign tb_data_input = 21795;
		#(CLK_PERIOD);
		assign tb_data_input = 21796;
		#(CLK_PERIOD);
		assign tb_data_input = 21797;
		#(CLK_PERIOD);
		assign tb_data_input = 21798;
		#(CLK_PERIOD);
		assign tb_data_input = 21799;
		#(CLK_PERIOD);
		assign tb_data_input = 21800;
		#(CLK_PERIOD);
		assign tb_data_input = 21801;
		#(CLK_PERIOD);
		assign tb_data_input = 21802;
		#(CLK_PERIOD);
		assign tb_data_input = 21803;
		#(CLK_PERIOD);
		assign tb_data_input = 21804;
		#(CLK_PERIOD);
		assign tb_data_input = 21805;
		#(CLK_PERIOD);
		assign tb_data_input = 21806;
		#(CLK_PERIOD);
		assign tb_data_input = 21807;
		#(CLK_PERIOD);
		assign tb_data_input = 21808;
		#(CLK_PERIOD);
		assign tb_data_input = 21809;
		#(CLK_PERIOD);
		assign tb_data_input = 21810;
		#(CLK_PERIOD);
		assign tb_data_input = 21811;
		#(CLK_PERIOD);
		assign tb_data_input = 21812;
		#(CLK_PERIOD);
		assign tb_data_input = 21813;
		#(CLK_PERIOD);
		assign tb_data_input = 21814;
		#(CLK_PERIOD);
		assign tb_data_input = 21815;
		#(CLK_PERIOD);
		assign tb_data_input = 21816;
		#(CLK_PERIOD);
		assign tb_data_input = 21817;
		#(CLK_PERIOD);
		assign tb_data_input = 21818;
		#(CLK_PERIOD);
		assign tb_data_input = 21819;
		#(CLK_PERIOD);
		assign tb_data_input = 21820;
		#(CLK_PERIOD);
		assign tb_data_input = 21821;
		#(CLK_PERIOD);
		assign tb_data_input = 21822;
		#(CLK_PERIOD);
		assign tb_data_input = 21823;
		#(CLK_PERIOD);
		assign tb_data_input = 21824;
		#(CLK_PERIOD);
		assign tb_data_input = 21825;
		#(CLK_PERIOD);
		assign tb_data_input = 21826;
		#(CLK_PERIOD);
		assign tb_data_input = 21827;
		#(CLK_PERIOD);
		assign tb_data_input = 21828;
		#(CLK_PERIOD);
		assign tb_data_input = 21829;
		#(CLK_PERIOD);
		assign tb_data_input = 21830;
		#(CLK_PERIOD);
		assign tb_data_input = 21831;
		#(CLK_PERIOD);
		assign tb_data_input = 21832;
		#(CLK_PERIOD);
		assign tb_data_input = 21833;
		#(CLK_PERIOD);
		assign tb_data_input = 21834;
		#(CLK_PERIOD);
		assign tb_data_input = 21835;
		#(CLK_PERIOD);
		assign tb_data_input = 21836;
		#(CLK_PERIOD);
		assign tb_data_input = 21837;
		#(CLK_PERIOD);
		assign tb_data_input = 21838;
		#(CLK_PERIOD);
		assign tb_data_input = 21839;
		#(CLK_PERIOD);
		assign tb_data_input = 21840;
		#(CLK_PERIOD);
		assign tb_data_input = 21841;
		#(CLK_PERIOD);
		assign tb_data_input = 21842;
		#(CLK_PERIOD);
		assign tb_data_input = 21843;
		#(CLK_PERIOD);
		assign tb_data_input = 21844;
		#(CLK_PERIOD);
		assign tb_data_input = 21845;
		#(CLK_PERIOD);
		assign tb_data_input = 21846;
		#(CLK_PERIOD);
		assign tb_data_input = 21847;
		#(CLK_PERIOD);
		assign tb_data_input = 21848;
		#(CLK_PERIOD);
		assign tb_data_input = 21849;
		#(CLK_PERIOD);


		if (tb_discrimination_parameter == 1'b0) begin
			$info("Test case 1 passed!");
		end else begin
			$info("Test case 1 failed, bro.");
		end

		#(2 * CLK_PERIOD); // Get away from time = 0.

		/* === Test Case 2 === 

		assign tb_useful_event_enable = 1'b1;
		assign tb_baseline_value = 12500;
		assign tb_current_maximum_value = 22500;

		#(CLK_PERIOD);

		if (tb_useful_event_out == 1'b1) begin
			$info("Test case 2 passed!");
		end else begin
			$info("Test case 2 failed, bro.");
		end

		#(2 * CLK_PERIOD); // Get away from time = 0.

		/* === Test Case 3 === 

		assign tb_useful_event_enable = 1'b1;
		assign tb_baseline_value = 12500;
		assign tb_current_maximum_value = 12000;

		#(CLK_PERIOD);

		if (tb_useful_event_out == 1'b0) begin
			$info("Test case 3 passed!");
		end else begin
			$info("Test case 3 failed, bro.");
		end

		#(2 * CLK_PERIOD); // Get away from time = 0.

		/* === Test Case 4 === 

		assign tb_tx_out = 1'b0;
		assign tb_sda_mode = 2'b11;

		#(CLK_PERIOD);

		if (tb_sda_out == tb_tx_out) begin
			$info("Test case 4 passed!");
		end else begin
			$info("Test case 4 failed, bro.");
		end

		#(2 * CLK_PERIOD); // Get away from time = 0. */

	end

endmodule
